`timescale 1ns / 1ps

`ifdef PRE_SYNTH_SIM
   `include "vsdbabysoc.v"
   `include "avsddac.v"
   `include "avsdpll.v"
   `include "rvmyth.v"
   `include "clk_gate.v"
`elsif POST_SYNTH_SIM
   `include "../../output/synth/vsdbabysoc.synth.v"
   `include "avsddac.v"
   `include "avsdpll.v"
   `include "../gls_model/primitives.v"
`else
   $error("Must define PRE_SYNTH_SIM or POST_SYNTH_SIM")
`endif

module vsdbabysoc_tb;
   reg       reset;
   reg       VCO_IN;
   reg       ENb_CP;
   reg       ENb_VCO;
   reg       REF;
   reg  real VREFL;
   reg  real VREFH;
   wire real OUT;

   vsdbabysoc uut (
      .OUT(OUT),
      .reset(reset),
      .VCO_IN(VCO_IN),
      .ENb_CP(ENb_CP),
      .ENb_VCO(ENb_VCO),
      .REF(REF),
      .VREFH(VREFH)
   );

   initial begin
      reset = 0;
      VREFL = 0.0;
      VREFH = 3.3;
      {REF, ENb_VCO, ENb_CP} = 0;
      VCO_IN = 1'b0;
      
      #20 reset = 1;
      #100 reset = 0;
      #10 ENb_CP = 1;
      #10 ENb_VCO = 1;
   end
   
   initial begin
`ifdef PRE_SYNTH_SIM
      $dumpfile("../../output/pre_synth_sim/pre_synth_sim.vcd");
`elsif POST_SYNTH_SIM
      $dumpfile("../../output/post_synth_sim/post_synth_sim.vcd");
`endif
      $dumpvars(0, vsdbabysoc_tb);
   end
 
   initial begin
      repeat(600) begin
         ENb_VCO = 1;
         #100 REF = ~REF;
         #(83.33/2) VCO_IN = ~VCO_IN;
      end
      $finish;
   end
   
endmodule
